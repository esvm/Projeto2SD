module PC(clk, out);

input wire clk;
output reg[3:0] out;

always @(posedge clk) begin
	if(out == 4'b1111) out = 4'b0000;
	else out = out + 1;
end

endmodule 