module registrador(In, cod, clk, out);
input[3:0] In;
input[1:0] cod;
input clk;
output[3:0] out;

endmodule
